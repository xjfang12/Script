`timescale 1ns/1ps
////////////////////////////////////////////////////////////////////////////////
//
// Filename:    test_tb.v
// Author:      FangXinjia
// Create Time: Mon Jul 15 13:32:24 2019
// Release:     First Release
// Project:     
// Modified:
//
//
//
// Description: 
//
//
//
//
////////////////////////////////////////////////////////////////////////////////
module test_tb; 
////////////////////////////////////////////////////////////////////////////////
// signal list
////////////////////////////////////////////////////////////////////////////////
reg        a;
reg        b;
reg        c;
reg        d;
reg  [3:0] e;
reg  [3:0] f;
reg  [3:0] g;
wire       h;
wire       i;
wire       j;
wire       l;
wire       m;
wire       n;
wire       o;
wire       p;
wire       q;


////////////////////////////////////////////////////////////////////////////////
// initial block
initial begin
  a = 0;
  b = 0;
  c = 0;
  d = 0;
  e = 0;
  f = 0;
  g = 0;
  #100;
end




////////////////////////////////////////////////////////////////////////////////
// UUT instance
////////////////////////////////////////////////////////////////////////////////
test u_test (
  .a(a),
  .b(b),
  .c(c),
  .d(d),
  .e(e),
  .f(f),
  .g(g),
  .h(h),
  .i(i),
  .j(j),
  .l(l),
  .m(m),
  .n(n),
  .o(o),
  .p(p),
  .q(q)
);



////////////////////////////////////////////////////////////////////////////////
// Clock Generate use if you need
////////////////////////////////////////////////////////////////////////////////
// always #5 clk = ~clk


endmodule
