`timescale 1ns/1ps
////////////////////////////////////////////////////////////////////////////////
//
// Filename:    test.v
// Author:      FangXinjia
// Create Time: Thu Mar 29 13:16:07 2018
// Release:     First Release
// Project:     
// Modified:
//
//
//
// Description: 
//
//
//
//
////////////////////////////////////////////////////////////////////////////////
module test (
	a,
	b,
	c,
	d,
	e, f, g,
	h,
	i,
	j,
	l,m,n,
	o,p,q

);

input a;
input b;
input c;
input d;
input [3:0] e,f,g;
output h;
output i;
output j;
output l,m,n;
inout o,p,q;

////////////////////////////////////////////////////////////////////////////////
// Local parameter define
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Wire and Reg define
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Main body
////////////////////////////////////////////////////////////////////////////////

endmodule
